module cla_tb;
reg [3:0] a;
reg [3:0] b;
reg c0;
wire [3:0] sum;
wire c_4;
cla uut(.sum(sum),.c_4(c_4),.a(a),.b(b),.c0(c0));
initial begin
a=0;
b=0;
c0=0;
#100;
a=1100;
b=0011;
c0=0;
end
endmodule
